../../axi4_lite_if.sv
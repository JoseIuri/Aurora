interface agentDummy_interface (input clock, reset);

    logic[8] in_data;
	logic[8] out_data;
	

    // modport port(
    // input   clock,
    // input   reset,
    // |-SIGNAL_NAME_PORT-|);

endinterface

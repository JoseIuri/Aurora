../../../axi4_types.sv